.include TSMC_180nm.txt
.param supply = 1.8

VCC net1 GND supply


*G0
MP9 o1 A0 net1 net1 CMOSP W=1.8u L=180nm
MP10 o1 B0 net1 net1 CMOSP W=1.8u L=180nm
MN9 o1 A0 o2 GND CMOSN W=0.9u L=180nm
MN10 o2 B0 GND GND CMOSN W=0.9u L=180nm
MP11 G0 o1 net1 net1 CMOSP W=1.8u L=180nm
MN11 G0 o1 GND GND CMOSN W=0.9u L=180nm

*G1
MP12 o3 A1 net1 net1 CMOSP W=1.8u L=180nm
MP13 o3 B1 net1 net1 CMOSP W=1.8u L=180nm
MN12 o3 A1 o4 GND CMOSN W=0.9u L=180nm
MN13 o4 B1 GND GND CMOSN W=0.9u L=180nm
MP14 G1 o3 net1 net1 CMOSP W=1.8u L=180nm
MN14 G1 o3 GND GND CMOSN W=0.9u L=180nm

*G2
MP15 o5 A2 net1 net1 CMOSP W=1.8u L=180nm
MP16 o5 B2 net1 net1 CMOSP W=1.8u L=180nm
MN15 o5 A2 o6 GND CMOSN W=0.9u L=180nm
MN16 o6 B2 GND GND CMOSN W=0.9u L=180nm
MP17 G2 o5 net1 net1 CMOSP W=1.8u L=180nm
MN17 G2 o5 GND GND CMOSN W=0.9u L=180nm

*G3
MP18 o7 A3 net1 net1 CMOSP W=1.8u L=180nm
MP19 o7 B3 net1 net1 CMOSP W=1.8u L=180nm
MN18 o7 A3 o8 GND CMOSN W=0.9u L=180nm
MN19 o8 B3 GND GND CMOSN W=0.9u L=180nm
MP20 G3 o7 net1 net1 CMOSP W=1.8u L=180nm
MN20 G3 o7 GND GND CMOSN W=0.9u L=180nm

*P0
MP21 o9 A0 net1 net1 CMOSP W=1.8u L=180nm
MN21 o9 A0 GND GND CMOSN W=0.9u L=180nm
MP22 P0 B0 A0 net1 CMOSP W=1.8u L=180nm
MN22 P0 B0 o9 GND CMOSN W=0.9u L=180nm
MP23 P0 A0 B0 net1 CMOSP W=1.8u L=180nm
MN23 B0 o9 P0 GND CMOSN W=0.9u L=180nm

*P1
MP24 o10 A1 net1 net1 CMOSP W=1.8u L=180nm
MN24 o10 A1 GND GND CMOSN W=0.9u L=180nm
MP25 P1 B1 A1 net1 CMOSP W=1.8u L=180nm
MN25 P1 B1 o10 GND CMOSN W=0.9u L=180nm
MP26 P1 A1 B1 net1 CMOSP W=1.8u L=180nm
MN26 B1 o10 P1 GND CMOSN W=0.9u L=180nm

*P2
MP27 o11 A2 net1 net1 CMOSP W=1.8u L=180nm
MN27 o11 A2 GND GND CMOSN W=0.9u L=180nm
MP28 P2 B2 A2 net1 CMOSP W=1.8u L=180nm
MN28 P2 B2 o11 GND CMOSN W=0.9u L=180nm
MP29 P2 A2 B2 net1 CMOSP W=1.8u L=180nm
MN29 B2 o11 P2 GND CMOSN W=0.9u L=180nm

*P3
MP30 o12 A3 net1 net1 CMOSP W=1.8u L=180nm
MN30 o12 A3 GND GND CMOSN W=0.9u L=180nm
MP31 P3 B3 A3 net1 CMOSP W=1.8u L=180nm
MN31 P3 B3 o12 GND CMOSN W=0.9u L=180nm
MP32 P3 A3 B3 net1 CMOSP W=1.8u L=180nm
MN32 B3 o12 P3 GND CMOSN W=0.9u L=180nm

*C1=G0+P0C0
MP33 o13 C0 net1 net1 CMOSP W=1.8u L=180nm
MP34 o13 P0 net1 net1 CMOSP W=1.8u L=180nm
MP35 o14 G0 o13 net1 CMOSP W=1.8u L=180nm
MN33 o14 P0 o15 GND CMOSN W=0.9u L=180nm
MN34 o15 C0 GND GND CMOSN W=0.9u L=180nm
MN35 o14 G0 GND GND CMOSN W=0.9u L=180nm
MP36 C1 o14 net1 net1 CMOSP W=1.8u L=180nm
MN36 C1 o14 GND GND CMOSN W=0.9u L=180nm

*C2=G1+P1C1=G1+P1(G0+POC0)
MP37 o16 P0 net1 net1 CMOSP W=1.8u L=180nm
MP38 o16 C0 net1 net1 CMOSP W=1.8u L=180nm
MP39 o17 G0 o16 net1 CMOSP W=1.8u L=180nm
MP40 o17 P1 net1 net1 CMOSP W=1.8u L=180nm
MP41 o18 G1 o17 net1 CMOSP W=1.8u L=180nm
MN37 o18 P1 o19 GND CMOSN W=0.9u L=180nm
MN38 019 P0 o20 GND CMOSN W=0.9u L=180nm
MN39 o20 C0 GND GND CMOSN W=0.9u L=180nm
MN40 o19 G0 GND GND CMOSN W=0.9u L=180nm
MN41 o18 G1 GND GND CMOSN W=0.9u L=180nm
MP42 C2 o18 net1 net1 CMOSP W=1.8u L=180nm
MN42 C2 o18 GND GND CMOSN W=0.9u L=180nm

*C3=G2+P2C2=G2+P2(G1+P1C1)=G2+P2[G1+P1(G0+P0C0)]
MP43 o21 P0 net1 net1 CMOSP W=1.8u L=180nm
MP44 o22 G0 o21 net1 CMOSP W=1.8u L=180nm
MP45 o23 G1 o22 net1 CMOSP W=1.8u L=180nm
MP46 o24 G2 o23 net1 CMOSP W=1.8u L=180nm
MP47 o21 C0 net1 net1 CMOSP W=1.8u L=180nm
MP48 o22 P1 net1 net1 CMOSP W=1.8u L=180nm
MP49 o23 P2 net1 net1 CMOSP W=1.8u L=180nm
MN43 o24 P2 o25 GND CMOSN W=0.9u L=180nm
MN44 o25 P1 o26 GND CMOSN W=0.9u L=180nm
MN45 o26 P0 o27 GND CMOSN W=0.9u L=180nm
MN46 o27 C0 GND GND CMOSN W=0.9u L=180nm
MN47 o26 G0 GND GND CMOSN W=0.9u L=180nm
MN48 o25 G1 GND GND CMOSN W=0.9u L=180nm
MN49 o24 G2 GND GND CMOSN W=0.9u L=180nm
MP50 C3 o24 net1 net1 CMOSP W=1.8u L=180nm
MN50 C3 o24 GND GND CMOSN W=0.9u L=180nm

*C4=G3+P3C3=G3+P3[G2+P2[G1+P1(G0+P0C0)]]
MP51 o28 P0 net1 net1 CMOSP W=1.8u L=180nm
MP52 o28 C0 net1 net1 CMOSP W=1.8u L=180nm
MP53 o29 G0 o28 net1 CMOSP W=1.8u L=180nm
MP54 o30 G1 o29 net1 CMOSP W=1.8u L=180nm
MP55 o31 G2 o30 net1 CMOSP W=1.8u L=180nm
MP56 o32 G3 o31 net1 CMOSP W=1.8u L=180nm
MP57 o29 P1 net1 net1 CMOSP W=1.8u L=180nm
MP58 o30 P2 net1 net1 CMOSP W=1.8u L=180nm
MP59 o31 P3 net1 net1 CMOSP W=1.8u L=180nm
MN51 o32 P3 o33 GND CMOSN W=0.9u L=180nm
MN52 o33 P2 o34 GND CMOSN W=0.9u L=180nm
MN53 o34 P1 o35 GND CMOSN W=0.9u L=180nm
MN54 o35 P0 o36 GND CMOSN W=0.9u L=180nm
MN55 o36 C0 GND GND CMOSN W=0.9u L=180nm
MN56 o32 G3 GND GND CMOSN W=0.9u L=180nm
MN57 o33 G2 GND GND CMOSN W=0.9u L=180nm
MN58 o34 G1 GND GND CMOSN W=0.9u L=180nm
MN59 o35 G0 GND GND CMOSN W=0.9u L=180nm
MP60 C4 o32 net1 net1 CMOSP W=1.8u L=180nm
MN60 C4 o32 GND GND CMOSN W=0.9u L=180nm



**S0=C0 XOR P0
MP61 o40 C0 net1 net1 CMOSP W=1.8u L=180nm
MN61 o40 C0 GND GND CMOSN W=0.9u L=180nm
MP62 S0 P0 C0 net1 CMOSP W=1.8u L=180nm
MN62 S0 P0 o40 GND CMOSN W=0.9u L=180nm
MP63 S0 C0 P0 net1 CMOSP W=1.8u L=180nm
MN63 P0 o40 S0 GND CMOSN W=0.9u L=180nm

**S1=C1 XOR P1
MP64 o41 C1 net1 net1 CMOSP W=1.8u L=180nm
MN64 o41 C1 GND GND CMOSN W=0.9u L=180nm
MP65 S1 P1 C1 net1 CMOSP W=1.8u L=180nm
MN65 S1 P1 o41 GND CMOSN W=0.9u L=180nm
MP66 S1 C1 P1 net1 CMOSP W=1.8u L=180nm
MN66 P1 o41 S1 GND CMOSN W=0.9u L=180nm

**S2=C2 XOR P2
MP67 o42 C2 net1 net1 CMOSP W=1.8u L=180nm
MN67 o42 C2 GND GND CMOSN W=0.9u L=180nm
MP68 S2 P2 C2 net1 CMOSP W=1.8u L=180nm
MN68 S2 P2 o42 GND CMOSN W=0.9u L=180nm
MP69 S2 C2 P2 net1 CMOSP W=1.8u L=180nm
MN69 P2 o42 S2 GND CMOSN W=0.9u L=180nm

**S3=C3 XOR P3
MP70 o43 C3 net1 net1 CMOSP W=1.8u L=180nm
MN70 o43 C3 GND GND CMOSN W=0.9u L=180nm
MP71 S3 P3 C3 net1 CMOSP W=1.8u L=180nm
MN71 S3 P3 o43 GND CMOSN W=0.9u L=180nm
MP72 S3 C3 P3 net1 CMOSP W=1.8u L=180nm
MN72 P3 o43 S3 GND CMOSN W=0.9u L=180nm

Vin1 A0 GND pulse(0 supply 0 1n 1n 0.1u 0.2u)
Vin2 B0 GND pulse(0 supply 0 1n 1n 0.2u 0.4u)
Vin3 A1 GND pulse(0 supply 0 1n 1n 0.1u 0.2u)
Vin4 B1 GND pulse(0 supply 0 1n 1n 0.2u 0.4u)
Vin5 A2 GND pulse(0 supply 0 1n 1n 0.1u 0.2u)
Vin6 B2 GND pulse(0 supply 0 1n 1n 0.2u 0.4u)
Vin7 A3 GND pulse(0 supply 0 1n 1n 0.1u 0.2u)
Vin8 B3 GND pulse(0 supply 0 1n 1n 0.2u 0.4u)
Vin9 C0 GND pulse (0 0 0 0.5p 0.5p 0.2u 0.4u)

Cap1 C1 GND 0.1p
Cap2 C2 GND 0.1p
Cap3 C3 GND 0.1p
Cap4 C4 GND 0.1p
Cap5 S0 GND 0.1p
Cap6 S1 GND 0.1p
Cap7 S2 GND 0.1p
Cap8 S3 GND 0.1p

.tran 1n 0.4u
.control
run

set curplottitle="Nanditha Merugu-2020102061"
plot v(C1)
set curplottitle="Nanditha Merugu-2020102061"
plot v(C2)
set curplottitle="Nanditha Merugu-2020102061"
plot v(C3)
set curplottitle="Nanditha Merugu-2020102061"
plot v(C4)
set curplottitle="Nanditha Merugu-2020102061"
plot v(S0)
set curplottitle="Nanditha Merugu-2020102061"
plot v(S1)
set curplottitle="Nanditha Merugu-2020102061"
plot v(S2)
set curplottitle="Nanditha Merugu-2020102061"
plot v(S3)
set curplottitle="Nanditha Merugu-2020102061"

.endc
.end








